magic
tech sky130A
timestamp 1725211376
<< nwell >>
rect -100 0 300 540
<< nmos >>
rect 95 -150 110 -50
<< pmos >>
rect 95 45 110 355
<< ndiff >>
rect 50 -60 95 -50
rect 50 -140 60 -60
rect 80 -140 95 -60
rect 50 -150 95 -140
rect 110 -60 155 -50
rect 110 -140 125 -60
rect 145 -140 155 -60
rect 110 -150 155 -140
<< pdiff >>
rect 45 345 95 355
rect 45 55 55 345
rect 80 55 95 345
rect 45 45 95 55
rect 110 345 160 355
rect 110 55 125 345
rect 150 55 160 345
rect 110 45 160 55
<< ndiffc >>
rect 60 -140 80 -60
rect 125 -140 145 -60
<< pdiffc >>
rect 55 55 80 345
rect 125 55 150 345
<< psubdiff >>
rect 40 -200 160 -185
rect 40 -230 55 -200
rect 145 -230 160 -200
rect 40 -245 160 -230
<< nsubdiff >>
rect 25 495 170 505
rect 25 445 45 495
rect 150 445 170 495
rect 25 435 170 445
<< psubdiffcont >>
rect 55 -230 145 -200
<< nsubdiffcont >>
rect 45 445 150 495
<< poly >>
rect 95 355 110 405
rect 95 10 110 45
rect 15 0 110 10
rect 15 -25 25 0
rect 50 -25 110 0
rect 15 -30 110 -25
rect 185 0 230 10
rect 185 -25 195 0
rect 220 -25 230 0
rect 185 -30 230 -25
rect 95 -50 110 -30
rect 95 -175 110 -150
<< polycont >>
rect 25 -25 50 0
rect 195 -25 220 0
<< locali >>
rect 25 495 170 505
rect 25 445 45 495
rect 150 445 170 495
rect 25 435 170 445
rect 45 345 90 435
rect 45 55 55 345
rect 80 55 90 345
rect 45 45 90 55
rect 115 345 160 355
rect 115 55 125 345
rect 150 55 160 345
rect 115 45 160 55
rect 15 0 60 10
rect 15 -25 25 0
rect 50 -25 60 0
rect 15 -30 60 -25
rect 120 -50 155 45
rect 185 0 230 10
rect 185 -25 195 0
rect 220 -25 230 0
rect 185 -30 230 -25
rect 50 -60 90 -50
rect 50 -140 60 -60
rect 80 -140 90 -60
rect 50 -185 90 -140
rect 115 -60 155 -50
rect 115 -140 125 -60
rect 145 -140 155 -60
rect 115 -150 155 -140
rect 50 -190 65 -185
rect 45 -200 65 -190
rect 110 -200 155 -190
rect 45 -230 55 -200
rect 145 -230 155 -200
rect 45 -235 65 -230
rect 110 -235 155 -230
rect 45 -240 155 -235
rect 50 -245 90 -240
<< viali >>
rect 60 445 105 495
rect 25 -25 50 0
rect 195 -25 220 0
rect 65 -200 110 -185
rect 65 -230 110 -200
rect 65 -235 110 -230
<< metal1 >>
rect -360 495 520 505
rect -360 445 60 495
rect 105 445 520 495
rect -360 435 520 445
rect -115 0 60 10
rect -115 -25 25 0
rect 50 -25 60 0
rect -115 -30 60 -25
rect 120 0 430 10
rect 120 -25 195 0
rect 220 -25 430 0
rect 120 -30 430 -25
rect -340 -185 540 -175
rect -340 -235 65 -185
rect 110 -235 540 -185
rect -340 -245 540 -235
<< labels >>
rlabel metal1 410 470 415 475 1 vdd
rlabel metal1 466 -220 500 -205 1 vcc
rlabel metal1 384 -15 418 0 1 out
<< end >>
